module hdmi_driver #(
    parameter N = 1
) ( 
    input sys_clk_i
);
    
endmodule