
module moduleName (
    
);
    
endmodule