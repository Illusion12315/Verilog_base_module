// ********************************************************************************** // 
//---------------------------------------------------------------------
// ������ת������ģ��
//---------------------------------------------------------------------
module bin2gray
#(
    parameter                           integer DATA_WIDTH = 256    
)
(
    input              [DATA_WIDTH-1:0] bin_i                      ,
    output             [DATA_WIDTH-1:0] gray_o                      
);

assign gray_o = (bin_i >> 1) ^ bin_i ;

endmodule